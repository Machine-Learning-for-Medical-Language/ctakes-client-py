ANAT|Anatomy|T024|Tissue
CHEM|Chemicals & Drugs|T195|Antibiotic