68235000|C0027424|Nasal congestion
64531003|C1260880|Rhinorrhea
49727002|C0010200|Coughing
11833005|C0850149|Dry Cough
28743005|C0239134|Productive Cough
62315008|C0011991|Diarrhea
84229001|C0015672|Fatigue
367391008|C0231218|Malaise
43724002|C0085593|Chills
43724002|C0036973|Shivering
103001002|C0687681|Feeling feverish
426000000|C1959900|Fever greater than 100.4 Fahrenheit
386661006|C0015967|Fever
274640006|C0085594|Chills and fever
25064002|C0018681|Headache
68962001|C0231528|Myalgia
82991003|C0281856|Myalgia
422587007|C0027497|Nausea
422400008|C0042963|Vomiting
16932000|C0027498|Nausea and vomiting
44169009|C0003126|Anosmia
36955009|C2364111|Ageusia
36955009|C0013378|Dysgeusia
267036007|C0013404|Dyspnea
162397003|C0242429|Sore throat