#CUI|TUI|CODE|SAB|STR|PREF
C0239134|T033|28743005|SNOMEDCT_US|Productive Cough|Cough
C0015672|T184|84229001|SNOMEDCT_US|Fatigue|Fatigue